package uart_package;

endpackage
