
interface serial_if;
  
    logic sdata;
    logic tick_rx;

endinterface: serial_if