
interface serial_if();

  logic sdata;
  logic handshake;
  logic tick_tx;
  logic tick_rx;

endinterface : serial_if
