module uart #(
    parameter SYSTEM_FREQUENCY = 100000000,
    parameter SAMPLING_RATE = 16
)(
    input clk,
    input reset_n,
    
    input [7:0] data_i,
    input tx_en_i,
    input rx_en_i,
    input start_tx_i,
    input [2:0] baud_sl_i,
    input  stop_bit_num,
    input [1:0] data_bit_num,
    input parity_en_i,
    input parity_type,
    
    // UART TX output
    output data_o,
    output data_o_valid
);

    // Internal signals
    logic tick_tx;
    logic tick_rx; 

    // Baud generator instance
    baud_generator #(
        .SYSTEM_FREQUENCY(SYSTEM_FREQUENCY),
        .SAMPLING_RATE(SAMPLING_RATE)
    ) baud_gen_inst (
        .clk(clk),
        .reset_n(reset_n),
        .baud_sl_i(baud_sl_i),
        .tick_tx(tick_tx),
        .tick_rx(tick_rx)
    );

    // UART transmitter instance
    wire tx;
    wire trans_fi_o;
    uart_transmitter uart_tx_inst (
        .clk(clk),
        .reset_n(reset_n),
        .start_tx_i(start_tx_i),
        .tx_en_i(tx_en_i),
        .parity_type_i(parity_type),
        .parity_en_i(parity_en_i),
        .data_i(data_i),
        .tick_i(tick_tx),
        .stop_bit_num_i(stop_bit_num),
        .data_bit_num_i(data_bit_num),
        .tx_o(tx),
        .trans_fi_o(trans_fi_o)
    );
    wire parity_err_o;
    wire stop_bit_err_o;
    uart_receiver inst_uart_receiver
        (
            .clk            (clk),
            .reset_n        (reset_n),
            .rx_en_i        (rx_en_i),
            .tick_i         (tick_rx),
            .parity_type_i  (parity_type),
            .parity_en_i    (parity_en_i),
            .tx_i           (tx),
            .stop_bit_num_i (stop_bit_num),
            .data_bit_num_i (data_bit_num),
            .data_o         (data_o),
            .data_o_valid   (data_o_valid),
            .parity_err_o   (parity_err_o),
            .stop_bit_err_o (stop_bit_err_o)
        );



endmodule
