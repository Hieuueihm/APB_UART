
interface serial_if;
  
    logic sdata;
    logic tick_rx;
    logic handshake;

endinterface: serial_if