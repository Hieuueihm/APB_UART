
interface serial_if();

  logic sdata;
  logic handshake;
  logic tick_tx;
  logic tick_rx;
  logic clk;
endinterface : serial_if
