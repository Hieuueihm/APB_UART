
interface serial_if;

  logic sdata;
  logic tick_rx;
  logic tick_tx;
  logic handshake;

endinterface : serial_if
