`define LOG(NAME, MSG) `uvm_info(NAME, MSG, UVM_LOW)
`define APB_AGENT_CFG "APB_AGENT_CFG"
`define APB_DRIVER     "APB_DRIVER"
`define APB_AGENT      "APB_AGENT"
`define APB_MONITOR    "APB_MONITOR"
`define APB_IF         "APB_INTERFACE"



`define UART_AGENT_CFG "UART_AGENT_CFG"
`define UART_DRIVER     "UART_DRIVER"
`define UART_AGENT      "UART_AGENT"
`define UART_MONITOR    "UART_MONITOR"


`define UART_ENV_CFG "UART_ENV_CFG"
`define UART_ENV      "UART_ENV"
`define UART_REG_CFG "UART_REG_CFG"
`define UART_REG      "UART_REG"

`define UART_TX_SCOREBOARD "UART_TX_SCOREBOARD"
`define UART_RX_SCOREBOARD "UART_RX_SCOREBOARD"