package uart_agent_pkg;
	
	import uvm_pkg::*;
	`include "uvm_macros.svh";
	// import common_def::*;

endpackage